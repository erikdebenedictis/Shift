  nRERL top level script
* [Under ngspice 36, { sS2, sQ2, snR, saa }.cir are an introduction to S2LAL, Q2LAL, and nRERL circuit.  Use files in vcs checked in h:mm PM d/mm/2022 (public)]

* Copyright 2022 Zettaflops, LLC

* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at

*     http://www.apache.org/licenses/LICENSE-2.0

* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* The top-level control is to switch which of the next lines are commented.
.param Ckt=4 T=27 Div=100 mn=1 mp=2                         $ defaults for control lines; nRERL does not benefit from a s-shaped ramp
.param o1=.15 h1=.15 o2=.30 h2=.30                          $ defaults for control lines; nRERL does not benefit from a s-shaped ramp
*.param      Vp=5v      MD=3        Vt=2.5v   Cg=1e-12    Cx=5e-18    wX=1        ww=60u      ll=.5u









*** RUN 1 Builtin BSIM 3
***param MD=3 J_S=1 Vp=9V       Hz=1e6      wX=1  ww=5u       ll=5u       Cw=.01p     Cb=5e-12    xl=9        xn=5  xh=5        yl=1e6      yn=1  yh=5e7
***param MD=5 Vt=.75v Vp=1.4v   Hz=1e6            wX=1  ww=500e-9   ll=150e-9   Cg=5e-15    Cx=5e-18    xl=.35       xn=1 xh=.35      yl=.4675    yn=-1 yh=.4675
*param MD=3 Vt=2.5v Vp=5.0v   Hz=1e6            wX=1  ww=500e-9   ll=150e-9   Cg=5e-13    Cx=5e-18    xl=5.0       xn=1 xh=5.0      yl=.4675    yn=-1 yh=.4675
* 0 Adia , 3 , 8.13859E-10 , 1.90592E-10 , 5 , 0.4675 , 5 , 0.25 , 5E-18 , 27 , 1 , 1 , 0.15 , 0.35 , 0.3 , 0.4675 , 31.607 4/16/22 7:09 4130
* 0 Adia , 3 , 5.35929E-10 , 1.31232E-10 , 5 , 0.4675 , 5 , 0.25 , 5E-18 , 27 , 1 , 1 , 0.15 , 0.15 , 0.3 , 0.3 , 31.21 4/18/22 5:38 4130

*** RUN 2 Speculative BSIM 4
***param MD=4 J_S=0 Vp=.275V    Hz=1e6      wX=1  ww=600e-9   ll=20e-9    Cw=.01p     Cb=5e-14    xl=.275     xn=5  xh=.175     yl=1e6      yn=1  yh=25e6
*param MD=4 Vt=.12v Vp=.40v   Hz=1e6            wX=1  ww=500e-9   ll=150e-9   Cg=5e-15    Cx=5e-18    xl=.35       xn=1 xh=.35      yl=.4675    yn=-1 yh=.4675
* 0 Adia , 4 , 5.60825E-14 , 3.41232E-14 , 0.4 , 0.4675 , 0.4 , 0.25 , 5E-18 , 27 , 1 , 1 , 0.15 , 0.35 , 0.3 , 0.4675 , 48.946 4/16/22 6:48 4130
* 0 Adia , 4 , 9.77748E-14 , 3.22176E-14 , 0.35 , 0.4675 , 0.35 , 0.25 , 5E-18 , 27 , 1 , 1 , 0.15 , 0.15 , 0.3 , 0.3 , 40.968 4/18/22 5:15 4130

*** RUN 3 Sky130 (this control line enabled by default)
.param MD=5 Vt=.75v Vp=2.8v   Hz=1e6            wX=1  ww=500e-9   ll=150e-9   Cg=5e-16    Cx=5e-17    xl=3.0      xn=3  xh=3.2      yl=.30      yn=-1 yh=.30
* 0 Adia , 5 , 5.87059E-13 , 3.1055E-14 , 3.1 , 0.3 , 3.1 , 0.25 , 5E-17 , 27 , 1 , 1 , 0.15 , 0.15 , 0.3 , 0.3 , 58.243 4/17/22 5:47 4130
* 1 Adia , 5 , 7.81334E-13 , 1.42033E-14 , 3.1 , 0.3 , 3.1 , 0.25 , 5E-17 , 27 , 1 , 1 , 0.15 , 0.15 , 0.3 , 0.3 , 94.7 4/18/22 5:13 4130







*** RUN 4 [undisclosed soi]
* Vtho on graph is .35 on scale of 1, but Vp = .8, so Vtho is .35*.8 = .28
*param MD=6 Vt=.28v Vp=0.8v   Hz=1e6            wX=1  ww=500e-9   ll=150e-9   Cg=2e-15    Cx=2e-16    xl=0.8       xn=1 xh=0.8      yl=.4675    yn=-1 yh=.4675
* 0 Adia , 6 , 6.60334E-14 , 1.16657E-14 , 0.8 , 0.4675 , 0.8 , 0.25 , 2E-16 , 27 , 1 , 1 , 0.15 , 0.15 , 0.3 , 0.3 , 120.101 4/17/22 3:54 4130
* 0 Adia , 6 , 9.29629E-14 , 1.30104E-14 , 0.8 , 0.4675 , 0.8 , 0.25 , 2E-16 , 27 , 1 , 1 , 0.15 , 0.15 , 0.3 , 0.3 , 109.089 4/18/22 5:24 4130



*PARAM MD=2 CKT=0 Vp=9.99V    Hz=1e4      T=27  wX=1  ww=5u       ll=5u       Cw=1e-17    Cb=100e-12  xl=9.99     xn=1  xh=9.99     yl=1e4      yn=1  yh=1e4

.param xvar=.15 yvar=.30                                    $ optional dummy variables that will be modified by the looping code in saa.cir
.param Vp=xvar $ h2=yvar

* The following equations are correct, but in the circuit Cg and Cx are in parallel with the simulated devices, which are not accounted for
.param b='Cg/(Cg+Cx)'                                       $ boosting factor [nRERL, between eq. (2) and eq. (3)]
.param m='Vp/Vt'                                            $ Vdd/Vt [nRERL, between Fig. 5 axis]
.param Vx='Vp*(1+b)-Vt'                                     $ Voltage of boost above Vdd [nRERL, between eq. (5)]
.param ACAP=0.001e-15                                       $ capacitive load on the data line

*** SUBCIRCUIT DEFINITIONS
* nRERL buffer [nRERL, Fig. 6a]
.SUBCKT nRERL f0 f1 f2 f3 X0P X0N X1P X1N nn1 nn2 nn3 nn4 GND PWR nsub psub ini='gg'
.ic V(nn1)='1.5*(vv-ini)' V(nn2)='1.5*vv'                   $ .ic V(a)={gg} V(a2)=ini
.ic V(nn4)='1.5*(vv-ini)' V(nn3)='1.5*vv'                   $ .ic V(a)={gg} V(a2)=ini
xM1  f1  X0P nn1 nsub nFET w=1 l=1                          $ logic switch
C01 X0P GND 'Cx'
C02 X0P f1 'Cg/2'
C03 X0P nn1 'Cg/2'
xM2  f1  X0N nn2 nsub nFET w=1 l=1                          $ logic switch
C11 X0N GND 'Cx'
C12 X0N f1 'Cg/2'
C13 X0N nn2 'Cg/2'
xM3  f2  X1P nn3 nsub nFET w=1 l=1                          $ logic switch
C21 X1P GND 'Cx'
C22 X1P f2 'Cg/2'
C23 X1P nn3 'Cg/2'
xM4  f2  X1N nn4 nsub nFET w=1 l=1                          $ logic switch
C31 X1N GND 'Cx'
C32 X1N f2 'Cg/2'
C33 X1N nn4 'Cg/2'
xM5  X1P f0  nn1 nsub nFET w=1 l=1                          $ isolation switch
xM6  X1N f0  nn2 nsub nFET w=1 l=1                          $ isolation switch
xM7  X0P f3  nn3 nsub nFET w=1 l=1                          $ isolation switch
xM8  X0N f3  nn4 nsub nFET w=1 l=1                          $ isolation switch
xM9  X1P X1N GND nsub nFET w=1 l=1                          $ clamp
xM10 X1N X1P GND nsub nFET w=1 l=1                          $ clamp
C40 X0P GND ACAP
C41 X0N GND ACAP
.ENDS nRERL

* A null nRERL buffer for implementing skips, [Complexity, Fig. 4ab]
.SUBCKT xRERL f0 f1 f2 f3 X0P X0N X1P X1N nn1 nn2 nn3 nn4 GND PWR nsub psub ini='gg'
r1 X0P X1P 0
r2 X0N X1N 0
.ENDS xRERL

.param va='gg'                                              $ initialization values for initialization to 1. Not sure these are right
.param vb='gg'
.param vc='gg'
.param vd='gg'
.param ve='gg'
.param vf='.67*vv'
.param vg='1.0*vv'
.param vh='1.0*vv'
.param vi='.67*vv'

*** TOP-LEVEL CIRCUIT
* for skips [complexity Fig. 4c] use a text editor to switch an nRERL to xRERL
x0  110 111 112 113 1000 2000 1001 2001 3001 3002 3003 3004 70 71 70 71 nRERL ini='va'
x1  111 112 113 114 1001 2001 1002 2002 3011 3012 3013 3014 70 71 70 71 nRERL ini='vb'
x2  112 113 114 115 1002 2002 1003 2003 3021 3022 3023 3024 70 71 70 71 nRERL ini='vc'
x3  113 114 115 116 1003 2003 1004 2004 3031 3032 3033 3034 70 71 70 71 nRERL ini='vd'
x4  114 115 116 117 1004 2004 1005 2005 3041 3042 3043 3044 70 71 70 71 nRERL ini='ve'
x5  115 116 117 110 1005 2005 1006 2006 3051 3052 3053 3054 70 71 70 71 nRERL ini='vf'
x6  116 117 110 111 1006 2006 1007 2007 3061 3062 3063 3064 70 71 70 71 nRERL ini='vg'
x7  117 110 111 112 1007 2007 1008 2008 3071 3072 3073 3074 70 71 70 71 nRERL ini='vh'

x8  110 111 112 113 1008 2008 1009 2009 3081 3082 3083 3084 70 71 70 71 nRERL ini='gg'
x9  111 112 113 114 1009 2009 1010 2010 3091 3092 3093 3094 70 71 70 71 nRERL ini='gg'
x10 112 113 114 115 1010 2010 1011 2011 3101 3102 3103 3104 70 71 70 71 nRERL ini='gg'
x11 113 114 115 116 1011 2011 1012 2012 3111 3112 3113 3114 70 71 70 71 nRERL ini='gg'
x12 114 115 116 117 1012 2012 1013 2013 3121 3122 3123 3124 70 71 70 71 nRERL ini='gg'
x13 115 116 117 110 1013 2013 1014 2014 3131 3132 3133 3134 70 71 70 71 nRERL ini='gg'
x14 116 117 110 111 1014 2014 1015 2015 3141 3142 3143 3144 70 71 70 71 nRERL ini='gg'
x15 117 110 111 112 1015 2015 1016 2016 3151 3152 3153 3154 70 71 70 71 nRERL ini='gg'

x16 110 111 112 113 1016 2016 1017 2017 3161 3162 3163 3164 70 71 70 71 nRERL ini='va'
x17 111 112 113 114 1017 2017 1018 2018 3171 3172 3173 3174 70 71 70 71 nRERL ini='vb'
x18 112 113 114 115 1018 2018 1019 2019 3181 3182 3183 3184 70 71 70 71 nRERL ini='vc'
x19 113 114 115 116 1019 2019 1020 2020 3191 3192 3193 3194 70 71 70 71 nRERL ini='vd'
x20 114 115 116 117 1020 2020 1021 2021 3201 3202 3203 3204 70 71 70 71 nRERL ini='ve'
x21 115 116 117 110 1021 2021 1022 2022 3211 3212 3213 3214 70 71 70 71 nRERL ini='vf'
x22 116 117 110 111 1022 2022 1023 2023 3221 3222 3223 3224 70 71 70 71 nRERL ini='vg'
x23 117 110 111 112 1023 2023 1000 2000 3231 3232 3233 3234 70 71 70 71 nRERL ini='vh'

r1000 1000 wv3_00 0
r1001 1001 wv3_01 0
r1002 1002 wv3_02 0
r1003 1003 wv3_03 0
r1004 1004 wv3_04 0
r1005 1005 wv3_05 0
r1006 1006 wv3_06 0
r1007 1007 wv3_07 0
r1008 1008 wv3_08 0
r1009 1009 wv3_09 0
r1010  110 wv3_10 0                                         $ the next 15 lines are a combination of 6-phase [nRERL, Fig 7] and 8-phase [Complexity]
r1011  111 wv3_11 0
r1012  112 wv3_12 0
r1013  113 wv3_13 0
r1014  114 wv3_14 0
r1015  115 wv3_15 0
r1016  116 wv3_16 0
r1017  117 wv3_17 0
r1018 1008 wv3_18 0
r1019 2008 wv3_19 0
r1020 1009 wv3_20 0
r1021 2009 wv3_21 0
r1022 3081 wv3_22 0
r1023 3083 wv3_23 0

r2000 2000 wv4_00 0
r2001 2001 wv4_01 0
r2002 2002 wv4_02 0
r2003 2003 wv4_03 0
r2004 2004 wv4_04 0
r2005 2005 wv4_05 0
r2006 2006 wv4_06 0
r2007 2007 wv4_07 0
r2008 3081 wv4_08 0
r2009 3082 wv4_09 0
r2010 3083 wv4_10 0
r2011 3084 wv4_11 0
r2012 3091 wv4_12 0
r2013 3092 wv4_13 0
r2014 3093 wv4_14 0
r2015 3094 wv4_15 0
r2016 3101 wv4_16 0
r2017 3102 wv4_17 0
r2018 3103 wv4_18 0
r2019 3104 wv4_19 0
r2020 3111 wv4_20 0
r2021 3112 wv4_21 0
r2022 3113 wv4_22 0
r2023 3114 wv4_23 0

* Cheapo initialization by overdriving some signals
.model switch1 sw vt=.1 ron=100k roff=1e12                     $ Ron and roff are repeating defaults. Seems to need the 1e12 value and e16 does not work
*s10 1000 124 123 70 switch1 on
*s11 2000 70 123 70 switch1 on
*s12 2008 124 123 70 switch1 on
*s13 1008 70 123 70 switch1 on
*s14 1016 124 123 70 switch1 on
*s15 2016 70 123 70 switch1 on

.inc saa.cir