* NGSPICE file created from qPhase11.ext - technology: sky130A

.subckt QAAmp11 S0T S0C S1T p1T Cl0 GN2 p0T p4T p2T Cl1 p3T p7T Vp T GND
X0 T S0C p1T GND sky130_fd_pr__nfet_01v8 ad=1.2025e+12p pd=9.8e+06u as=3.75e+11p ps=2.6e+06u w=450000u l=150000u
X1 GND Cl0 T GND sky130_fd_pr__nfet_01v8 ad=5.025e+11p pd=4.2e+06u as=0p ps=0u w=450000u l=150000u
X2 S1T p0T T GND sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=0p ps=0u w=450000u l=150000u
X3 T S0T GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X4 S1T p4T T Vp sky130_fd_pr__pfet_01v8 ad=2.25e+11p pd=1.9e+06u as=2.7e+11p ps=2.1e+06u w=450000u l=150000u
X5 T S0T p1T Vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.25e+11p ps=1.9e+06u w=450000u l=150000u
C0 GN2 p0T 0.10fF
C1 Vp p1T 0.36fF
C2 S0C p1T 0.08fF
C3 p1T T 0.41fF
C4 p2T p1T 0.08fF
C5 Cl0 p1T 0.15fF
C6 p3T p7T 0.17fF
C7 S0T p1T 0.62fF
C8 Vp p7T 0.01fF
C9 S1T Vp 0.06fF
C10 S1T p4T 0.17fF
C11 Vp p4T 0.11fF
C12 p7T T 0.04fF
C13 S1T Cl1 0.04fF
C14 S0C p3T 0.06fF
C15 S1T T 0.16fF
C16 p4T Cl1 0.43fF
C17 Cl0 p7T 0.50fF
C18 Vp T 0.09fF
C19 S1T GN2 0.04fF
C20 S0T p7T 0.04fF
C21 p4T T 0.14fF
C22 Cl0 p3T 0.53fF
C23 Vp GN2 0.12fF
C24 Vp p2T 0.20fF
C25 S0T p3T 0.04fF
C26 p4T GN2 0.35fF
C27 p4T p2T 0.16fF
C28 Cl1 T 0.04fF
C29 S0C T 0.02fF
C30 S0T Vp 0.26fF
C31 GN2 Cl1 0.14fF
C32 p2T Cl1 0.07fF
C33 S0T p4T 0.02fF
C34 GN2 T 0.04fF
C35 p2T T 0.06fF
C36 S1T p0T 0.25fF
C37 Cl0 S0C 0.01fF
C38 Cl0 T 0.11fF
C39 GN2 p2T 0.19fF
C40 S0T S0C 0.04fF
C41 S0T T 0.09fF
C42 p4T p0T 0.22fF
C43 Cl1 p0T 0.48fF
C44 p7T p1T 0.14fF
C45 S0T Cl0 0.18fF
C46 p3T p1T 0.05fF
C47 S1T p1T 0.01fF
C48 Cl1 GND 0.19fF
C49 GN2 GND 0.16fF
C50 p2T GND 0.15fF
C51 p7T GND 0.47fF
C52 p3T GND 0.25fF
C53 S1T GND 0.42fF
C54 p1T GND 0.68fF
C55 p0T GND 0.44fF
C56 p4T GND 0.44fF
C57 S0T GND 0.71fF
C58 S0C GND 0.30fF
C59 Cl0 GND 0.61fF
C60 Vp GND 0.58fF
C61 T GND 0.61fF
.ends

.subckt qLatch11 AT AC QT QC p0T p1T p7T GN2 PWR p2T p3T p4T GND Cl0 Cl1
XQAAmp11_0 AC AT QC p1T Cl0 GN2 p0T p4T p2T Cl1 p3T p7T PWR QAAmp11_0/T GND QAAmp11
XQAAmp11_1 AT AC QT p1T Cl0 GN2 p0T p4T p2T Cl1 p3T p7T PWR QAAmp11_1/T GND QAAmp11
C0 AT p1T 0.09fF
C1 AT AC 0.36fF
C2 QT QC 0.02fF
C3 AC p1T 0.03fF
C4 QAAmp11_0/T QAAmp11_1/T 0.31fF
C5 AT QAAmp11_0/T 0.05fF
C6 QAAmp11_1/T QC 0.01fF
C7 AT QAAmp11_1/T 0.01fF
C8 QAAmp11_0/T p1T 0.07fF
C9 p1T QAAmp11_1/T 0.07fF
C10 QAAmp11_0/T QT 0.01fF
C11 AC QAAmp11_1/T 0.05fF
C12 QT GND 0.45fF
C13 AT GND 1.27fF
C14 AC GND 1.45fF
C15 PWR GND 1.40fF
C16 QAAmp11_1/T GND 0.61fF
C17 Cl1 GND 0.36fF
C18 GN2 GND 0.31fF
C19 p2T GND 0.29fF
C20 p7T GND 0.93fF
C21 p3T GND 0.49fF
C22 QC GND 0.45fF
C23 p1T GND 1.35fF
C24 p0T GND 0.88fF
C25 p4T GND 0.87fF
C26 Cl0 GND 1.21fF
C27 QAAmp11_0/T GND 0.61fF
.ends

.subckt qPhase11 S0T S0C S1T S1C p0T p0C p1T Cl1 p2T Cl2 p3T p3C GN2 PWR
XqLatch11_0 S0T S0C S1T S1C p0T p1T p3C GN2 PWR p2T p3T p0C GN2 Cl1 Cl2 qLatch11
XqLatch11_1 S1T S1C S0T S0C p3T p2T p0C GN2 PWR p1T p0T p3C GN2 Cl2 Cl1 qLatch11
C0 S0T S0C 0.67fF
C1 S1T S1C 0.18fF
C2 Cl1 S0T 0.20fF
C3 S0T p3C 0.14fF
C4 Cl2 S1C 0.02fF
C5 S0T p1T 0.04fF
C6 Cl1 S0C 0.14fF
C7 S1T p0T 0.20fF
C8 p2T S1C 0.06fF
C9 S0T p3T 0.26fF
C10 S0C p3T 0.19fF
C11 Cl2 S1T 0.15fF
C12 S0T GN2 2.20fF
C13 S1T GN2 2.41fF
C14 S1C GN2 2.66fF
C15 qLatch11_1/QAAmp11_1/T GN2 0.61fF
C16 qLatch11_1/QAAmp11_0/T GN2 0.61fF
C17 S0C GN2 2.44fF
C18 PWR GN2 3.19fF
C19 qLatch11_0/QAAmp11_1/T GN2 0.61fF
C20 Cl2 GN2 1.55fF
C21 p2T GN2 1.59fF
C22 p3C GN2 1.79fF
C23 p3T GN2 1.36fF
C24 p1T GN2 1.63fF
C25 p0T GN2 1.33fF
C26 p0C GN2 1.79fF
C27 Cl1 GN2 1.57fF
C28 qLatch11_0/QAAmp11_0/T GN2 0.61fF
.ends

